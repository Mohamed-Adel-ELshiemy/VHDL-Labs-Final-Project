 -- Import the necessary packages
LIBRARY ieee;
USE std.textio.ALL;
use ieee.std_logic_textio.all;
USE ieee.numeric_bit.ALL;
USE ieee.std_logic_1164.ALL;
-- uSE WORK.pack_a.ALL;


entity NBitMultiplierDivider_TB is
end entity NBitMultiplierDivider_TB;

architecture tb_arch of NBitMultiplierDivider_TB is
  constant N : positive := 8; -- Number of bits

  signal a       : std_logic_vector(N-1 downto 0);
  signal b       : std_logic_vector(N-1 downto 0);
  signal op      : std_logic;
  signal m       : std_logic_vector(2*N-1 downto 0); -- Update the size to accommodate the larger result
  signal r       : std_logic_vector(N-1 downto 0);
  signal error   : std_logic;
  signal busy    : std_logic;
  signal valid   : std_logic;
  
  -- Clock process
  constant CLK_PERIOD : time := 10 ns;
  signal clk : std_logic := '0';

-- Declare a line variable for writing results
signal result_line : line;

begin

  DUT: entity work.NBitMultiplierDivider
    generic map (
      N => N
    )
    port map (
      a     => a,
      b     => b,
      op    => op,
      m     => m,
      r     => r,
      error => error,
      busy  => busy,
      valid => valid
    );

  -- Clock process
  clk_process: process
  begin
    while now < 1000 ns loop
      clk <= '0';
      wait for CLK_PERIOD/2;
      clk <= '1';
      wait for CLK_PERIOD/2;
    end loop;
    wait;
  end process clk_process;

  -- Stimulus process
  stimulus_process: process
  begin
    -- Initialize inputs
    a <= (others => '0');
    b <= (others => '0');
    op <= '0';
    wait for CLK_PERIOD;

    -- Test multiplication
    a <= (others => '0'); -- Example operand values
    b <= (others => '0');
    a(N-1 downto N/2) <= "1101"; -- Update specific bits for test case
    b(N-1 downto N/2) <= "1010";
    op <= '0';
    wait for CLK_PERIOD;
    
    -- Test division
    a <= (others => '0'); -- Example operand values
    b <= (others => '0');
    a(N-1 downto N/2) <= "10101"; -- Update specific bits for test case
    b(N-1 downto N/2) <= "0110";
    op <= '1';
    wait for CLK_PERIOD;

    -- Additional test cases...

    wait;
  end process stimulus_process;

-- Monitor process
monitor_process: process
  variable result_line : line;
begin
  while true loop
    wait until valid = '1';
    
    -- Clear the line variable
    textio.reset(result_line);
    
    -- Write the results to the line variable
    write(result_line, "Result: m = ");
    write(result_line, to_string(unsigned(m)));
    write(result_line, ", r = ");
    write(result_line, to_string(unsigned(r)));
    
    -- Report the result line
    report "Result: " & to_string(result_line);
    
    wait;
  end loop;
end process monitor_process;

end architecture tb_arch;